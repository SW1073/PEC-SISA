LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;

PACKAGE package_tlb IS

    CONSTANT W_SEL_VIRTUAL      : std_logic := '0';
    CONSTANT W_SEL_PHYSICAL     : std_logic := '1';

END package_tlb;

PACKAGE BODY package_tlb IS

END package_tlb;


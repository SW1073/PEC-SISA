LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;        --Esta libreria sera necesaria si usais conversiones TO_INTEGER
USE ieee.std_logic_unsigned.ALL; --Esta libreria sera necesaria si usais conversiones CONV_INTEGER
USE work.package_io.ALL;

ENTITY controladores_IO IS
    PORT (
        boot       : IN  STD_LOGIC;
        CLOCK_50   : IN  STD_LOGIC;
        addr_io    : IN  STD_LOGIC_VECTOR(7  DOWNTO 0);
        wr_io      : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
        rd_io      : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        wr_out     : IN  STD_LOGIC;
        rd_in      : IN  STD_LOGIC;
        SW         : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        KEY        : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        hex        : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        hex_on     : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        led_verdes : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        led_rojos  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        ps2_clk    : inout STD_LOGIC;
        ps2_data   : inout STD_LOGIC);
END controladores_IO;

ARCHITECTURE Structure OF controladores_IO IS

    COMPONENT keyboard_controller is
        Port (clk        : in    STD_LOGIC;
              reset      : in    STD_LOGIC;
              ps2_clk    : inout STD_LOGIC;
              ps2_data   : inout STD_LOGIC;
              read_char  : out   STD_LOGIC_VECTOR (7 downto 0);
              clear_char : in    STD_LOGIC;
              data_ready : out   STD_LOGIC);
    end COMPONENT;

    TYPE Mat IS ARRAY (255 DOWNTO 0) OF std_logic_vector(15 DOWNTO 0);
    SIGNAL registers : Mat := (OTHERS => (OTHERS => '0'));

    SIGNAL s_ps2_ascii_code : std_logic_vector(7 downto 0);
    SIGNAL s_ps2_clear_char : std_logic;
    SIGNAL s_ps2_data_ready : std_logic;

    SIGNAL contador_ciclos          : std_logic_vector(15 downto 0);
    SIGNAL contador_milisegundos    : std_logic_vector(15 downto 0);
BEGIN

    process(CLOCK_50)
    begin
        if rising_edge(CLOCK_50) then
            if contador_ciclos=0 then
                contador_ciclos<=x"C350"; -- tiempo de ciclo=20ns(50Mhz) 1ms=50000ciclos
                if contador_milisegundos>0 then
                    contador_milisegundos <= contador_milisegundos-1;
                end if;
            else
                contador_ciclos <= contador_ciclos-1;
            end if;
        end if;
    end process;

    PROCESS (CLOCK_50) IS
    BEGIN
        IF rising_edge(CLOCK_50) THEN
            registers(PORT_KEY)(3 downto 0) <= KEY(3 DOWNTO 0);
            registers(PORT_SW)(7 downto 0) <= SW(7 DOWNTO 0);
            registers(PORT_RAND) <= contador_ciclos;
            registers(PORT_TIMER) <= contador_milisegundos;

            IF wr_out = '1' AND addr_io /= PORT_KEY AND addr_io /= PORT_SW THEN
                if addr_io = PORT_PS2_DATA_VALID THEN
                    registers(conv_integer(addr_io)) <= x"0000";
                    s_ps2_clear_char <= '0';
                ELSE
                    registers(conv_integer(addr_io)) <= wr_io;
                END IF;
            END IF;

            IF s_ps2_data_ready = '1' THEN
                registers(PORT_PS2_DATA)(7 downto 0) <= s_ps2_ascii_code;
                registers(PORT_PS2_DATA_VALID) <= x"FFFF";
                s_ps2_clear_char <= '1';
            END IF;
        END IF;
    END PROCESS;

    -- Read con enable
    rd_io <= registers(conv_integer(addr_io)) WHEN rd_in = '1' ELSE x"0000";

    hex <= registers(PORT_HEX)(15 downto 0);
    hex_on <= registers(PORT_HEX_OFF)(3 downto 0);
    led_verdes <= registers(PORT_GREEN_LEDS)(7 downto 0);
    led_rojos <= registers(PORT_RED_LEDS)(7 downto 0);



    keyboard_controller0: keyboard_controller PORT MAP(
        clk         => CLOCK_50,
        reset       => boot,
        ps2_clk     => ps2_clk,
        ps2_data    => ps2_data,
        read_char   => s_ps2_ascii_code,
        clear_char  => s_ps2_clear_char,
        data_ready  => s_ps2_data_ready
    );

END Structure;
